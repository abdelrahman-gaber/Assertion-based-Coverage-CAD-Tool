library verilog;
use verilog.vl_types.all;
entity bind_assertions is
end bind_assertions;
