library verilog;
use verilog.vl_types.all;
entity Coverage is
    port(
        clkw            : in     vl_logic;
        clksd           : in     vl_logic
    );
end Coverage;
